//
// File: hvl_standard_vip.sv
//
// Generated from Mentor VIP Configurator (20230807)
// Generated using Mentor VIP Library ( 2023.3_1 : 08/18/2023:20:00 )
//
module hvl_standard_vip;
    import uvm_pkg::*;
    
    `include "test_packages.svh"
    
    initial
    begin
        run_test();
    end

endmodule: hvl_standard_vip
