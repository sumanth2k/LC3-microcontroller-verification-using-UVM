//
// File: test_packages.svh
//
// Generated from Mentor VIP Configurator (20230807)
// Generated using Mentor VIP Library ( 2023.3_1 : 08/18/2023:20:00 )
//

import standard_vip_pkg::*;

// Add other packages here as required
