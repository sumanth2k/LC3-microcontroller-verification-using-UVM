//
// File: standard_vip_pkg.sv
//
// Generated from Mentor VIP Configurator (20230807)
// Generated using Mentor VIP Library ( 2023.3_1 : 08/18/2023:20:00 )
//
package standard_vip_pkg;
    import uvm_pkg::*;
    
    `include "uvm_macros.svh"
    
    import addr_map_pkg::*;
    
    import standard_vip_params_pkg::*;
    import mvc_pkg::*;
    import mgc_axi4_v1_0_pkg::*;
    
    `include "standard_vip_env_config.svh"
    `include "standard_vip_env.svh"
    `include "standard_vip_vseq_base.svh"
    `include "standard_vip_test_base.svh"
endpackage: standard_vip_pkg
